//////////////////////////////////////////////
// Project Name:     DDFS verilog
//                   
// Group:            
// Author(s):        Francesco Urbani
// 
// Create Date:      Mon Jan 14 18:09:39 W. Europe Daylight Time 2019
// Design Name: 
// Module Name:      lut_clk
// Target Devices:   Intel MAX10 10M50DAF484C7G
// Tool versions: 
// Description:      
//
// THIS FILE IS AUTOGENERATED BY LUT_generator.py
// WARNING! All changes made in this file might be lost!
//
// Revision:
//////////////////////////////////////////////


module lut_clk
#(
    parameter      N = 17,
    parameter      M = 1
)
(
    input wire   [N-1:0]     lut_line,
    output reg   [M-1:0]     lut_data
);
    

always @ (*) 
begin

    lut_data = (lut_line < 2**(N-1) ? 1 : 0);
    
end
endmodule
    