---------------------------------------------
-- Title       : LUT_DDFS_SG_4096x6
-- Project     : DDFS
---------------------------------------------
-- File        : LUT_DDFS_SG_4096x6.vhd
-- Language    : VHDL
-- Author(s)   : francescourbani
-- Company     : 
-- Created     : Wed May 16 20:11:47 CEST 2018
---------------------------------------------
-- Description : LUT for DDFS
--        N_FW : 12
--       lines : 4096
--        N_YQ : 6
--       SG_UN : SG
--         lsb : 0.03225806451612903
---------------------------------------------


-- new LUT with 1/4 of the full elements

library ieee;
use ieee.std_logic_1164.all;
-- use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;



entity Q_LUT is
	port (
		LUT_line : in  std_logic_vector(11 downto 0);
		LUT_data : out std_logic_vector(5 downto 0) 
	);
end Q_LUT;

architecture rtl of Q_LUT is
	type LUT_t is array (natural range 0 to 1023) of integer;
	constant LUT: LUT_t := (
		0 => 0,
		1 => 0,
		2 => 0,
		3 => 0,
		4 => 0,
		5 => 0,
		6 => 0,
		7 => 0,
		8 => 0,
		9 => 0,
		10 => 0,
		11 => 0,
		12 => 0,
		13 => 0,
		14 => 0,
		15 => 0,
		16 => 0,
		17 => 0,
		18 => 0,
		19 => 0,
		20 => 0,
		21 => 0,
		22 => 1,
		23 => 1,
		24 => 1,
		25 => 1,
		26 => 1,
		27 => 1,
		28 => 1,
		29 => 1,
		30 => 1,
		31 => 1,
		32 => 1,
		33 => 1,
		34 => 1,
		35 => 1,
		36 => 1,
		37 => 1,
		38 => 1,
		39 => 1,
		40 => 1,
		41 => 1,
		42 => 1,
		43 => 2,
		44 => 2,
		45 => 2,
		46 => 2,
		47 => 2,
		48 => 2,
		49 => 2,
		50 => 2,
		51 => 2,
		52 => 2,
		53 => 2,
		54 => 2,
		55 => 2,
		56 => 2,
		57 => 2,
		58 => 2,
		59 => 2,
		60 => 2,
		61 => 2,
		62 => 2,
		63 => 2,
		64 => 3,
		65 => 3,
		66 => 3,
		67 => 3,
		68 => 3,
		69 => 3,
		70 => 3,
		71 => 3,
		72 => 3,
		73 => 3,
		74 => 3,
		75 => 3,
		76 => 3,
		77 => 3,
		78 => 3,
		79 => 3,
		80 => 3,
		81 => 3,
		82 => 3,
		83 => 3,
		84 => 3,
		85 => 4,
		86 => 4,
		87 => 4,
		88 => 4,
		89 => 4,
		90 => 4,
		91 => 4,
		92 => 4,
		93 => 4,
		94 => 4,
		95 => 4,
		96 => 4,
		97 => 4,
		98 => 4,
		99 => 4,
		100 => 4,
		101 => 4,
		102 => 4,
		103 => 4,
		104 => 4,
		105 => 4,
		106 => 5,
		107 => 5,
		108 => 5,
		109 => 5,
		110 => 5,
		111 => 5,
		112 => 5,
		113 => 5,
		114 => 5,
		115 => 5,
		116 => 5,
		117 => 5,
		118 => 5,
		119 => 5,
		120 => 5,
		121 => 5,
		122 => 5,
		123 => 5,
		124 => 5,
		125 => 5,
		126 => 5,
		127 => 6,
		128 => 6,
		129 => 6,
		130 => 6,
		131 => 6,
		132 => 6,
		133 => 6,
		134 => 6,
		135 => 6,
		136 => 6,
		137 => 6,
		138 => 6,
		139 => 6,
		140 => 6,
		141 => 6,
		142 => 6,
		143 => 6,
		144 => 6,
		145 => 6,
		146 => 6,
		147 => 6,
		148 => 6,
		149 => 7,
		150 => 7,
		151 => 7,
		152 => 7,
		153 => 7,
		154 => 7,
		155 => 7,
		156 => 7,
		157 => 7,
		158 => 7,
		159 => 7,
		160 => 7,
		161 => 7,
		162 => 7,
		163 => 7,
		164 => 7,
		165 => 7,
		166 => 7,
		167 => 7,
		168 => 7,
		169 => 7,
		170 => 7,
		171 => 8,
		172 => 8,
		173 => 8,
		174 => 8,
		175 => 8,
		176 => 8,
		177 => 8,
		178 => 8,
		179 => 8,
		180 => 8,
		181 => 8,
		182 => 8,
		183 => 8,
		184 => 8,
		185 => 8,
		186 => 8,
		187 => 8,
		188 => 8,
		189 => 8,
		190 => 8,
		191 => 8,
		192 => 8,
		193 => 9,
		194 => 9,
		195 => 9,
		196 => 9,
		197 => 9,
		198 => 9,
		199 => 9,
		200 => 9,
		201 => 9,
		202 => 9,
		203 => 9,
		204 => 9,
		205 => 9,
		206 => 9,
		207 => 9,
		208 => 9,
		209 => 9,
		210 => 9,
		211 => 9,
		212 => 9,
		213 => 9,
		214 => 9,
		215 => 10,
		216 => 10,
		217 => 10,
		218 => 10,
		219 => 10,
		220 => 10,
		221 => 10,
		222 => 10,
		223 => 10,
		224 => 10,
		225 => 10,
		226 => 10,
		227 => 10,
		228 => 10,
		229 => 10,
		230 => 10,
		231 => 10,
		232 => 10,
		233 => 10,
		234 => 10,
		235 => 10,
		236 => 10,
		237 => 11,
		238 => 11,
		239 => 11,
		240 => 11,
		241 => 11,
		242 => 11,
		243 => 11,
		244 => 11,
		245 => 11,
		246 => 11,
		247 => 11,
		248 => 11,
		249 => 11,
		250 => 11,
		251 => 11,
		252 => 11,
		253 => 11,
		254 => 11,
		255 => 11,
		256 => 11,
		257 => 11,
		258 => 11,
		259 => 11,
		260 => 12,
		261 => 12,
		262 => 12,
		263 => 12,
		264 => 12,
		265 => 12,
		266 => 12,
		267 => 12,
		268 => 12,
		269 => 12,
		270 => 12,
		271 => 12,
		272 => 12,
		273 => 12,
		274 => 12,
		275 => 12,
		276 => 12,
		277 => 12,
		278 => 12,
		279 => 12,
		280 => 12,
		281 => 12,
		282 => 12,
		283 => 13,
		284 => 13,
		285 => 13,
		286 => 13,
		287 => 13,
		288 => 13,
		289 => 13,
		290 => 13,
		291 => 13,
		292 => 13,
		293 => 13,
		294 => 13,
		295 => 13,
		296 => 13,
		297 => 13,
		298 => 13,
		299 => 13,
		300 => 13,
		301 => 13,
		302 => 13,
		303 => 13,
		304 => 13,
		305 => 13,
		306 => 14,
		307 => 14,
		308 => 14,
		309 => 14,
		310 => 14,
		311 => 14,
		312 => 14,
		313 => 14,
		314 => 14,
		315 => 14,
		316 => 14,
		317 => 14,
		318 => 14,
		319 => 14,
		320 => 14,
		321 => 14,
		322 => 14,
		323 => 14,
		324 => 14,
		325 => 14,
		326 => 14,
		327 => 14,
		328 => 14,
		329 => 14,
		330 => 15,
		331 => 15,
		332 => 15,
		333 => 15,
		334 => 15,
		335 => 15,
		336 => 15,
		337 => 15,
		338 => 15,
		339 => 15,
		340 => 15,
		341 => 15,
		342 => 15,
		343 => 15,
		344 => 15,
		345 => 15,
		346 => 15,
		347 => 15,
		348 => 15,
		349 => 15,
		350 => 15,
		351 => 15,
		352 => 15,
		353 => 15,
		354 => 16,
		355 => 16,
		356 => 16,
		357 => 16,
		358 => 16,
		359 => 16,
		360 => 16,
		361 => 16,
		362 => 16,
		363 => 16,
		364 => 16,
		365 => 16,
		366 => 16,
		367 => 16,
		368 => 16,
		369 => 16,
		370 => 16,
		371 => 16,
		372 => 16,
		373 => 16,
		374 => 16,
		375 => 16,
		376 => 16,
		377 => 16,
		378 => 16,
		379 => 17,
		380 => 17,
		381 => 17,
		382 => 17,
		383 => 17,
		384 => 17,
		385 => 17,
		386 => 17,
		387 => 17,
		388 => 17,
		389 => 17,
		390 => 17,
		391 => 17,
		392 => 17,
		393 => 17,
		394 => 17,
		395 => 17,
		396 => 17,
		397 => 17,
		398 => 17,
		399 => 17,
		400 => 17,
		401 => 17,
		402 => 17,
		403 => 17,
		404 => 18,
		405 => 18,
		406 => 18,
		407 => 18,
		408 => 18,
		409 => 18,
		410 => 18,
		411 => 18,
		412 => 18,
		413 => 18,
		414 => 18,
		415 => 18,
		416 => 18,
		417 => 18,
		418 => 18,
		419 => 18,
		420 => 18,
		421 => 18,
		422 => 18,
		423 => 18,
		424 => 18,
		425 => 18,
		426 => 18,
		427 => 18,
		428 => 18,
		429 => 18,
		430 => 18,
		431 => 19,
		432 => 19,
		433 => 19,
		434 => 19,
		435 => 19,
		436 => 19,
		437 => 19,
		438 => 19,
		439 => 19,
		440 => 19,
		441 => 19,
		442 => 19,
		443 => 19,
		444 => 19,
		445 => 19,
		446 => 19,
		447 => 19,
		448 => 19,
		449 => 19,
		450 => 19,
		451 => 19,
		452 => 19,
		453 => 19,
		454 => 19,
		455 => 19,
		456 => 19,
		457 => 19,
		458 => 20,
		459 => 20,
		460 => 20,
		461 => 20,
		462 => 20,
		463 => 20,
		464 => 20,
		465 => 20,
		466 => 20,
		467 => 20,
		468 => 20,
		469 => 20,
		470 => 20,
		471 => 20,
		472 => 20,
		473 => 20,
		474 => 20,
		475 => 20,
		476 => 20,
		477 => 20,
		478 => 20,
		479 => 20,
		480 => 20,
		481 => 20,
		482 => 20,
		483 => 20,
		484 => 20,
		485 => 20,
		486 => 21,
		487 => 21,
		488 => 21,
		489 => 21,
		490 => 21,
		491 => 21,
		492 => 21,
		493 => 21,
		494 => 21,
		495 => 21,
		496 => 21,
		497 => 21,
		498 => 21,
		499 => 21,
		500 => 21,
		501 => 21,
		502 => 21,
		503 => 21,
		504 => 21,
		505 => 21,
		506 => 21,
		507 => 21,
		508 => 21,
		509 => 21,
		510 => 21,
		511 => 21,
		512 => 21,
		513 => 21,
		514 => 21,
		515 => 22,
		516 => 22,
		517 => 22,
		518 => 22,
		519 => 22,
		520 => 22,
		521 => 22,
		522 => 22,
		523 => 22,
		524 => 22,
		525 => 22,
		526 => 22,
		527 => 22,
		528 => 22,
		529 => 22,
		530 => 22,
		531 => 22,
		532 => 22,
		533 => 22,
		534 => 22,
		535 => 22,
		536 => 22,
		537 => 22,
		538 => 22,
		539 => 22,
		540 => 22,
		541 => 22,
		542 => 22,
		543 => 22,
		544 => 22,
		545 => 23,
		546 => 23,
		547 => 23,
		548 => 23,
		549 => 23,
		550 => 23,
		551 => 23,
		552 => 23,
		553 => 23,
		554 => 23,
		555 => 23,
		556 => 23,
		557 => 23,
		558 => 23,
		559 => 23,
		560 => 23,
		561 => 23,
		562 => 23,
		563 => 23,
		564 => 23,
		565 => 23,
		566 => 23,
		567 => 23,
		568 => 23,
		569 => 23,
		570 => 23,
		571 => 23,
		572 => 23,
		573 => 23,
		574 => 23,
		575 => 23,
		576 => 23,
		577 => 23,
		578 => 24,
		579 => 24,
		580 => 24,
		581 => 24,
		582 => 24,
		583 => 24,
		584 => 24,
		585 => 24,
		586 => 24,
		587 => 24,
		588 => 24,
		589 => 24,
		590 => 24,
		591 => 24,
		592 => 24,
		593 => 24,
		594 => 24,
		595 => 24,
		596 => 24,
		597 => 24,
		598 => 24,
		599 => 24,
		600 => 24,
		601 => 24,
		602 => 24,
		603 => 24,
		604 => 24,
		605 => 24,
		606 => 24,
		607 => 24,
		608 => 24,
		609 => 24,
		610 => 24,
		611 => 24,
		612 => 25,
		613 => 25,
		614 => 25,
		615 => 25,
		616 => 25,
		617 => 25,
		618 => 25,
		619 => 25,
		620 => 25,
		621 => 25,
		622 => 25,
		623 => 25,
		624 => 25,
		625 => 25,
		626 => 25,
		627 => 25,
		628 => 25,
		629 => 25,
		630 => 25,
		631 => 25,
		632 => 25,
		633 => 25,
		634 => 25,
		635 => 25,
		636 => 25,
		637 => 25,
		638 => 25,
		639 => 25,
		640 => 25,
		641 => 25,
		642 => 25,
		643 => 25,
		644 => 25,
		645 => 25,
		646 => 25,
		647 => 25,
		648 => 25,
		649 => 26,
		650 => 26,
		651 => 26,
		652 => 26,
		653 => 26,
		654 => 26,
		655 => 26,
		656 => 26,
		657 => 26,
		658 => 26,
		659 => 26,
		660 => 26,
		661 => 26,
		662 => 26,
		663 => 26,
		664 => 26,
		665 => 26,
		666 => 26,
		667 => 26,
		668 => 26,
		669 => 26,
		670 => 26,
		671 => 26,
		672 => 26,
		673 => 26,
		674 => 26,
		675 => 26,
		676 => 26,
		677 => 26,
		678 => 26,
		679 => 26,
		680 => 26,
		681 => 26,
		682 => 26,
		683 => 26,
		684 => 26,
		685 => 26,
		686 => 26,
		687 => 26,
		688 => 26,
		689 => 26,
		690 => 27,
		691 => 27,
		692 => 27,
		693 => 27,
		694 => 27,
		695 => 27,
		696 => 27,
		697 => 27,
		698 => 27,
		699 => 27,
		700 => 27,
		701 => 27,
		702 => 27,
		703 => 27,
		704 => 27,
		705 => 27,
		706 => 27,
		707 => 27,
		708 => 27,
		709 => 27,
		710 => 27,
		711 => 27,
		712 => 27,
		713 => 27,
		714 => 27,
		715 => 27,
		716 => 27,
		717 => 27,
		718 => 27,
		719 => 27,
		720 => 27,
		721 => 27,
		722 => 27,
		723 => 27,
		724 => 27,
		725 => 27,
		726 => 27,
		727 => 27,
		728 => 27,
		729 => 27,
		730 => 27,
		731 => 27,
		732 => 27,
		733 => 27,
		734 => 27,
		735 => 28,
		736 => 28,
		737 => 28,
		738 => 28,
		739 => 28,
		740 => 28,
		741 => 28,
		742 => 28,
		743 => 28,
		744 => 28,
		745 => 28,
		746 => 28,
		747 => 28,
		748 => 28,
		749 => 28,
		750 => 28,
		751 => 28,
		752 => 28,
		753 => 28,
		754 => 28,
		755 => 28,
		756 => 28,
		757 => 28,
		758 => 28,
		759 => 28,
		760 => 28,
		761 => 28,
		762 => 28,
		763 => 28,
		764 => 28,
		765 => 28,
		766 => 28,
		767 => 28,
		768 => 28,
		769 => 28,
		770 => 28,
		771 => 28,
		772 => 28,
		773 => 28,
		774 => 28,
		775 => 28,
		776 => 28,
		777 => 28,
		778 => 28,
		779 => 28,
		780 => 28,
		781 => 28,
		782 => 28,
		783 => 28,
		784 => 28,
		785 => 28,
		786 => 28,
		787 => 28,
		788 => 28,
		789 => 29,
		790 => 29,
		791 => 29,
		792 => 29,
		793 => 29,
		794 => 29,
		795 => 29,
		796 => 29,
		797 => 29,
		798 => 29,
		799 => 29,
		800 => 29,
		801 => 29,
		802 => 29,
		803 => 29,
		804 => 29,
		805 => 29,
		806 => 29,
		807 => 29,
		808 => 29,
		809 => 29,
		810 => 29,
		811 => 29,
		812 => 29,
		813 => 29,
		814 => 29,
		815 => 29,
		816 => 29,
		817 => 29,
		818 => 29,
		819 => 29,
		820 => 29,
		821 => 29,
		822 => 29,
		823 => 29,
		824 => 29,
		825 => 29,
		826 => 29,
		827 => 29,
		828 => 29,
		829 => 29,
		830 => 29,
		831 => 29,
		832 => 29,
		833 => 29,
		834 => 29,
		835 => 29,
		836 => 29,
		837 => 29,
		838 => 29,
		839 => 29,
		840 => 29,
		841 => 29,
		842 => 29,
		843 => 29,
		844 => 29,
		845 => 29,
		846 => 29,
		847 => 29,
		848 => 29,
		849 => 29,
		850 => 29,
		851 => 29,
		852 => 29,
		853 => 29,
		854 => 29,
		855 => 29,
		856 => 29,
		857 => 29,
		858 => 30,
		859 => 30,
		860 => 30,
		861 => 30,
		862 => 30,
		863 => 30,
		864 => 30,
		865 => 30,
		866 => 30,
		867 => 30,
		868 => 30,
		869 => 30,
		870 => 30,
		871 => 30,
		872 => 30,
		873 => 30,
		874 => 30,
		875 => 30,
		876 => 30,
		877 => 30,
		878 => 30,
		879 => 30,
		880 => 30,
		881 => 30,
		882 => 30,
		883 => 30,
		884 => 30,
		885 => 30,
		886 => 30,
		887 => 30,
		888 => 30,
		889 => 30,
		890 => 30,
		891 => 30,
		892 => 30,
		893 => 30,
		894 => 30,
		895 => 30,
		896 => 30,
		897 => 30,
		898 => 30,
		899 => 30,
		900 => 30,
		901 => 30,
		902 => 30,
		903 => 30,
		904 => 30,
		905 => 30,
		906 => 30,
		907 => 30,
		908 => 30,
		909 => 30,
		910 => 30,
		911 => 30,
		912 => 30,
		913 => 30,
		914 => 30,
		915 => 30,
		916 => 30,
		917 => 30,
		918 => 30,
		919 => 30,
		920 => 30,
		921 => 30,
		922 => 30,
		923 => 30,
		924 => 30,
		925 => 30,
		926 => 30,
		927 => 30,
		928 => 30,
		929 => 30,
		930 => 30,
		931 => 30,
		932 => 30,
		933 => 30,
		934 => 30,
		935 => 30,
		936 => 30,
		937 => 30,
		938 => 30,
		939 => 30,
		940 => 30,
		941 => 30,
		942 => 30,
		943 => 30,
		944 => 30,
		945 => 30,
		946 => 30,
		947 => 30,
		948 => 30,
		949 => 30,
		950 => 30,
		951 => 30,
		952 => 30,
		953 => 30,
		954 => 30,
		955 => 30,
		956 => 30,
		957 => 30,
		958 => 30,
		959 => 30,
		960 => 30,
		961 => 30,
		962 => 30,
		963 => 30,
		964 => 30,
		965 => 30,
		966 => 30,
		967 => 30,
		968 => 30,
		969 => 30,
		970 => 30,
		971 => 30,
		972 => 30,
		973 => 30,
		974 => 30,
		975 => 30,
		976 => 30,
		977 => 30,
		978 => 30,
		979 => 30,
		980 => 30,
		981 => 30,
		982 => 30,
		983 => 30,
		984 => 30,
		985 => 30,
		986 => 30,
		987 => 30,
		988 => 30,
		989 => 30,
		990 => 30,
		991 => 30,
		992 => 30,
		993 => 30,
		994 => 30,
		995 => 30,
		996 => 30,
		997 => 30,
		998 => 30,
		999 => 30,
		1000 => 30,
		1001 => 30,
		1002 => 30,
		1003 => 30,
		1004 => 30,
		1005 => 30,
		1006 => 30,
		1007 => 30,
		1008 => 30,
		1009 => 30,
		1010 => 30,
		1011 => 30,
		1012 => 30,
		1013 => 30,
		1014 => 30,
		1015 => 30,
		1016 => 30,
		1017 => 30,
		1018 => 30,
		1019 => 30,
		1020 => 30,
		1021 => 30,
		1022 => 30,
		1023 => 30
);

begin
	LUT_data <= std_logic_vector(TO_SIGNED(LUT(TO_INTEGER(unsigned(LUT_line))), 6));
end rtl;
